module Decoder_5to32(S,m);
	input[4:0]S;
	output[32:0]m;

	//00000// 
	assign m[0] = ~S[4] & ~S[3] & ~S[2] & ~S[1] & ~S[0];
	//00001// 
	assign m[1] = ~S[4] & ~S[3] & ~S[2] & ~S[1] & S[0];
	//00010// 
	assign m[2] = ~S[4] & ~S[3] & ~S[2] & S[1] & ~S[0];
	//00011// 
	assign m[3] = ~S[4] & ~S[3] & ~S[2] & S[1] & S[0];
	//00100// 
	assign m[4] = ~S[4] & ~S[3] & S[2] & ~S[1] & ~S[0];
	//00101// 
	assign m[5] = ~S[4] & ~S[3] & S[2] & ~S[1] & S[0];
	//00110// 
	assign m[6] = ~S[4] & ~S[3] & S[2] & S[1] & ~S[0];
	//00111// 
	assign m[7] = ~S[4] & ~S[3] & S[2] & S[1] & S[0];
	//01000// 
	assign m[8] = ~S[4] & S[3] & ~S[2] & ~S[1] & ~S[0];
	//01001// 
	assign m[9] = ~S[4] & S[3] & ~S[2] & ~S[1] & S[0];
	//01010// 
	assign m[10] = ~S[4] & S[3] & ~S[2] & S[1] & ~S[0];
	//01011// 
	assign m[11] = ~S[4] & S[3] & ~S[2] & S[1] & S[0];
	//01100// 
	assign m[12] = ~S[4] & S[3] & S[2] & ~S[1] & ~S[0];
	//01101//
	assign m[13] = ~S[4] & S[3] & S[2] & ~S[1] & S[0];
	//01110// 
	assign m[14] = ~S[4] & S[3] & S[2] & S[1] & ~S[0];
	//01111// 
	assign m[15] = ~S[4] & S[3] & S[2] & S[1] & S[0];
	//10000// 
	assign m[16] = S[4] & ~S[3] & ~S[2] & ~S[1] & ~S[0];
	//10001// 
	assign m[17] = S[4] & ~S[3] & ~S[2] & ~S[1] & S[0];
	//10010// 
	assign m[18] = S[4] & ~S[3] & ~S[2] & S[1] & ~S[0];
	//10011// 
	assign m[19] = S[4] & ~S[3] & ~S[2] & S[1] & S[0];
	//10100//
	assign m[20] = S[4] & ~S[3] & S[2] & ~S[1] & ~S[0];
	//10101// 
	assign m[21] = S[4] & ~S[3] & S[2] & ~S[1] & S[0];
	//10110//
	assign m[22] = S[4] & ~S[3] & S[2] & S[1] & ~S[0];
	//10111//
	assign m[23] = S[4] & ~S[3] & S[2] & S[1] & S[0];
	//11000// 
	assign m[24] = S[4] & S[3] & ~S[2] & ~S[1] & ~S[0];
	//11001// 
	assign m[25] = S[4] & S[3] & ~S[2] & ~S[1] & S[0];
	//11010// 
	assign m[26] = S[4] & S[3] & ~S[2] & S[1] & ~S[0];
	//11011// 
	assign m[27] = S[4] & S[3] & ~S[2] & S[1] & S[0];
	//11100//
	assign m[28] = S[4] & S[3] & S[2] & ~S[1] & ~S[0];
	//11101// 
	assign m[29] = S[4] & S[3] & S[2] & ~S[1] & S[0];
	//11110// 
	assign m[30] = S[4] & S[3] & S[2] & S[1] & ~S[0];
	//11111// 
	assign m[31] = S[4] & S[3] & S[2] & S[1] & S[0];
endmodule