module Mux_32to1(X,S,Y);
	input[31:0] X;
	input[4:0] S;
	output reg Y;

always@(X or S)
	begin
		case (S)
			5'b00000: Y <= X[0];
			5'b00001: Y <= X[1];
			5'b00010: Y <= X[2];
			5'b00011: Y <= X[3];
			5'b00100: Y <= X[4];
			5'b00101: Y <= X[5];
			5'b00110: Y <= X[6];
			5'b00111: Y <= X[7];
			
			5'b01000: Y <= X[8];
			5'b01001: Y <= X[9];
			5'b01010: Y <= X[10];
			5'b01011: Y <= X[11];
			5'b01100: Y <= X[12];
			5'b01101: Y <= X[13];
			5'b01110: Y <= X[14];
			5'b01111: Y <= X[15];
			
			5'b10000: Y <= X[16];
			5'b10001: Y <= X[17];
			5'b10010: Y <= X[18];
			5'b10011: Y <= X[19];
			5'b10100: Y <= X[20];
			5'b10101: Y <= X[21];
			5'b10110: Y <= X[22];
			5'b10111: Y <= X[23];
			
			5'b11000: Y <= X[24];
			5'b11001: Y <= X[25];
			5'b11010: Y <= X[26];
			5'b11011: Y <= X[27];
			5'b11100: Y <= X[28];
			5'b11101: Y <= X[29];
			5'b11110: Y <= X[30];
			5'b11111: Y <= X[31];
			

		endcase
	end
endmodule
